library IEEE;  
use IEEE.STD_LOGIC_1164.all; 
use IEEE.STD_LOGIC_UNSIGNED.all;

entity AUTOMAT is
	port (CLK, START, SEL_MODE, USA, BUTON_AUTO, BUTON_TEMPERATURA, BUTON_VITEZA, PRESPALARE_MANUAL, CLATIRE_SUPL_MANUAL: in STD_LOGIC;
	TEMPERATURA, VITEZA: inout INTEGER;	
	PRESPALARE, CLATIRE_SUPL, USA_BLOCATA: inout STD_LOGIC;  
	TIMP_TOTAL: inout NATURAL;
	ACTIV: out STD_LOGIC;
	ROTIRE, ALIMENTARE, INCALZIRE, EVACUARE, PRESPALARE_OUT, CLATIRE_SUPL_OUT: out STD_LOGIC;
	A_TO_G: out STD_LOGIC_VECTOR(6 downto 0);
	AN: out STD_LOGIC_VECTOR(3 downto 0));
end AUTOMAT;

architecture AUTOMAT_ARCH of AUTOMAT is	

--constante timpi
constant TIMP_SPALARE_PRINCIPALA: INTEGER := 120;
constant TIMP_CLATIRE: INTEGER := 60;
constant TIMP_CENTRIFUGARE: INTEGER := 60;
constant TIMP_PRESPALARE: INTEGER := 60;
constant TIMP_APA: INTEGER := 6;  

--divizor
component CLOCK_DIVIDER
	port (MCLK, CLR: in STD_LOGIC;
	CLK_DIVIZAT, CLK_DIVIZAT_AFIS: out STD_LOGIC);
end component; 	 

--clock-uri divizate
signal CLK_DIV: STD_LOGIC; 
signal CLK_DIV_AF: STD_LOGIC;
 
--debounce
component DEBOUNCE4_PUSH_BUTTONS
	port (CCLK, CLR: in STD_LOGIC; --clk divizat
	INP: in STD_LOGIC; 
	OUTP: out STD_LOGIC);
end component;		

--semnalele corecte de la butoane (debounced)
signal BUTON_AUTO_D, BUTON_TEMPERATURA_D, BUTON_VITEZA_D, START_D: STD_LOGIC;

--preluare date input
component GET_DATA
	port (MODE, BUTON_P, BUTON_T, BUTON_V, PRESPALARE_MANUAL, CLATIRE_MANUAL: in STD_LOGIC;
	PRESPALARE, CLATIRE_SUPL: out STD_LOGIC;
	VITEZA, TEMPERATURA: out INTEGER);
end component;	   

--calculare timp total 
component TIME_CALC
	port (TEMPERATURA, TIMP_SPALARE_PRINCIPALA, TIMP_CLATIRE, TIMP_CENTRIFUGARE, TIMP_PRESPALARE, TIMP_APA: in INTEGER;
	PRESPALARE, CLATIRE_SUPL: in STD_LOGIC;
	TIMP: out NATURAL);
end component;

--logica de stari
component NEXT_STATE_LOGIC
	port(START, PRESPALARE, CLATIRE_SUPL, USA, CLK: in STD_LOGIC; 
	TEMPERATURA: in INTEGER;
	PRESPALARE_OUT, CLATIRE_SUPL_OUT, ACTIV, ROTIRE, ALIMENTARE, INCALZIRE, EVACUARE, USA_BLOCATA: out STD_LOGIC);
end component; 

--timer
component TIMP_AFISOR
	port(CLK, START, USA: in STD_LOGIC;
	TIMP_IN: in NATURAL;
	TIMP_NATURAL: out NATURAL;
	TIMP: out STD_LOGIC_VECTOR(11 downto 0));	
end component;

--afisor
component AFISOR
	port (CLK: in STD_LOGIC;	   
	TIMP: in NATURAL;
	UNITATI, ZECI, SUTE, MII: in STD_LOGIC_VECTOR(3 downto 0);
	A_TO_G: out STD_LOGIC_VECTOR(6 downto 0);
	AN: out STD_LOGIC_VECTOR(3 downto 0));
end component; 

--conversia
component BIN_TO_BCD is
	port(BINAR: in STD_LOGIC_VECTOR(11 downto 0);
	UNITATI: out STD_LOGIC_VECTOR(3 downto 0);
	ZECI: out STD_LOGIC_VECTOR(3 downto 0);
	SUTE: out STD_LOGIC_VECTOR(3 downto 0);	
	MII: out STD_LOGIC_VECTOR(3 downto 0));
end component;

signal TIMP_AFIS: STD_LOGIC_VECTOR(11 downto 0);
signal TIMP_NATURAL: NATURAL;
signal UNITATI, ZECI, SUTE, MII: STD_LOGIC_VECTOR(3 downto 0);

begin  

DIVIZARE_CLK: CLOCK_DIVIDER port map (CLK, '0', CLK_DIV, CLK_DIV_AF); 
DEBOUNCE_AUTO: DEBOUNCE4_PUSH_BUTTONS port map (CLK_DIV, '0', BUTON_AUTO, BUTON_AUTO_D);
DEBOUNCE_TEMPERATURA: DEBOUNCE4_PUSH_BUTTONS port map (CLK_DIV, '0', BUTON_TEMPERATURA, BUTON_TEMPERATURA_D);
DEBOUNCE_VITEZA: DEBOUNCE4_PUSH_BUTTONS port map (CLK_DIV, '0', BUTON_VITEZA, BUTON_VITEZA_D);	
DEBOUNCE_START: DEBOUNCE4_PUSH_BUTTONS port map (CLK_DIV, '0', START, START_D);	
GET_INPUT: GET_DATA port map (SEL_MODE, BUTON_AUTO_D, BUTON_TEMPERATURA_D, BUTON_VITEZA_D, PRESPALARE_MANUAL, CLATIRE_SUPL_MANUAL, PRESPALARE, CLATIRE_SUPL, VITEZA, TEMPERATURA);
CALC_TIMP: TIME_CALC port map (TEMPERATURA, TIMP_SPALARE_PRINCIPALA, TIMP_CLATIRE, TIMP_CENTRIFUGARE, TIMP_PRESPALARE, TIMP_APA, PRESPALARE, CLATIRE_SUPL, TIMP_TOTAL);
STARE_NXT: NEXT_STATE_LOGIC port map (START_D, PRESPALARE, CLATIRE_SUPL, USA, CLK_DIV, TEMPERATURA, PRESPALARE_OUT, CLATIRE_SUPL_OUT, ACTIV, ROTIRE, ALIMENTARE, INCALZIRE, EVACUARE, USA_BLOCATA); 
TIMER: TIMP_AFISOR port map (CLK_DIV, START_D, USA, TIMP_TOTAL, TIMP_NATURAL, TIMP_AFIS);
AFISOR_7SEGM: AFISOR port map (CLK_DIV_AF, TIMP_NATURAL, UNITATI, ZECI, SUTE, MII, A_TO_G, AN);	
COMP: BIN_TO_BCD port map (TIMP_AFIS, UNITATI, ZECI, SUTE, MII);

end AUTOMAT_ARCH;